module power_pack2 #(parameter WIDTH=20,
										 HEIGHT=20, 
										 box_size = 7'd64) 
	 (input wire 			clk,
	  input wire 			reset,
	  input wire			eaten,
	  input wire			spawn,
	  input wire [10:0]	hcount,
	  input wire [9:0]	vcount,
	  input wire [10:0]	randx,
	  input wire [9:0]	randy,
	  output reg [10:0]	rx,
	  output reg [9:0]	ry,
	  output reg [9:0]	r2pixel,
	  output reg [1:0]	mode,
	  output wire			randop
	  );
	 
	reg			display;
	wire			x_valid, y_valid;
	reg randop_reg;  
	reg [7:0] color;
	wire [7:0] randnum;
	
	parameter SHRINK	= 	2'b00;
	parameter BOOST	= 	2'b01;
	parameter idk		= 	2'b10;
	parameter SHIELD	=	2'b11; 	
	
	
	parameter COLOR_SHRINK	= 	8'b000_000_11;
	parameter COLOR_BOOST	=	8'b000_101_10;
	parameter COLOR_IDK		=	8'b111_000_11;
	parameter COLOR_SHIELD	=	8'b111_100_00;
	
	
	randgen pptype_gen(.clk(clk), .LFSR(randnum));
	  
	always @(posedge clk)
		begin
			if(reset || (spawn && !eaten)) begin
				mode <= randnum[1:0];
				//mode <= SHIELD;
				case(mode)
					SHRINK: begin
						color <= COLOR_SHRINK;
						end
					BOOST: begin
						color <= COLOR_BOOST;
						end
					SHIELD: begin
						color <= COLOR_SHIELD;
						end
					idk: begin
						color <= COLOR_IDK;
						end
					endcase
				display <= 1;
				rx <= randx;//700;
				ry <= randy;//500;
				randop_reg <= 1;
				end
			else if(eaten) begin
				//display <= 0;
				rx <= 0;
				ry <= 0;
				end
			else
				randop_reg <= 0;
			end
	  
	always @(hcount or vcount) 
		begin
			if ((hcount >= rx && hcount < (rx+WIDTH)) && (vcount >= ry && vcount < (ry+HEIGHT))) begin
				if(display)
					r2pixel = color;
				else
					r2pixel = 0;
				end
			else 
				r2pixel= 0;	
			end
			
	assign randop = randop_reg;
	
endmodule


module shield(
	input wire clk,
	input wire reset,
	input wire active,
	input wire [10:0] hcount, paddle_x,
	input wire [9:0]  vcount, paddle_y,
	input wire [9:0] paddle_width, paddle_height,
	output reg [7:0] pixel
	);

	reg [10:0] rx, height;
	reg [9:0]  ry, width;

	parameter COLOR = 8'b111_100_00;
	parameter BORDER = 10;
	
	always @(posedge clk)
		begin
			rx <= 100;//paddle_x;
			ry <= 100;//paddle_y;
			width <= 50;//paddle_width;
			height <= 50;//paddle_height;
			end			

	always @(hcount or vcount) 
		begin
			if(active) begin
				//if((hcount >= rx - BORDER) && hcount < rx && (vcount >= ry - BORDER) && (vcount < ry + height + BORDER)) begin
				//if ((hcount >= (rx - 4'd10) && hcount < rx) && ((vcount >= ry - 4'd10) && vcount < (ry + height + 4'd10))) begin
				if ((hcount >= 90 && hcount < 110) && (vcount >= 90 && vcount < 160)) begin
					pixel = COLOR;
					end
				end
			else pixel = 0;
			end
	
endmodule
